LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY C_60_H IS
    PORT(
		CLK		:IN std_logic;
		DIN1: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		DIN0: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        CLK_60	:OUT std_logic);
END;

ARCHITECTURE BH OF C_60_H IS
SIGNAL	clk_out:	STD_LOGIC;
SIGNAL	M1,M0,S1,S0:	STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	M1 <= DIN1(7 DOWNTO 4);
	M0 <= DIN1(3 DOWNTO 0);
	S1<=DIN0(7 DOWNTO 4);
	S0<=DIN0(3 DOWNTO 0);
	PROCESS(clk)
	BEGIN
		IF (CLK'EVENT AND clk='1') THEN
			IF (M1=5 AND M0=9 AND S1=5 AND S0=9) THEN
				clk_out <= '1';
			ELSE CLK_OUT<='0';
			END IF;
		END IF;
	END PROCESS;
	clk_60 <= clk_out;
END BH;