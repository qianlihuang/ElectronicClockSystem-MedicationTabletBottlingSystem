LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TWO_FOUR IS
	PORT(SETTIME0,SETTIME1,SETTIME_EN:IN STD_LOGIC;
		Y0,Y1,Y2,Y3:OUT STD_LOGIC);
END TWO_FOUR;

ARCHITECTURE BH OF TWO_FOUR IS
BEGIN
	PROCESS(SETTIME_EN,SETTIME1,SETTIME0)
	BEGIN
		IF(SETTIME1='0' AND SETTIME0='0' AND SETTIME_EN='1')THEN
			Y3<='1';
			Y2<='1';
			Y1<='1';
			Y0<='0';
		ELSIF(SETTIME1='0' AND SETTIME0='1' AND SETTIME_EN='1')THEN
			Y3<='1';
			Y2<='1';
			Y1<='0';
			Y0<='1';
		ELSIF(SETTIME1='1' AND SETTIME0='0' AND SETTIME_EN='1')THEN
			Y3<='1';
			Y2<='0';
			Y1<='1';
			Y0<='1';
		ELSIF(SETTIME1='1' AND SETTIME0='1' AND SETTIME_EN='1')THEN
			Y3<='0';
			Y2<='1';
			Y1<='1';
			Y0<='1';
		ELSE
			Y3<='1';
			Y2<='1';
			Y1<='1';
			Y0<='1';
		END IF;
	END PROCESS;
END BH;