LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY C_60 IS
    PORT(
		CLK		:IN std_logic;
		DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        CLK_60	:OUT std_logic);
END;

ARCHITECTURE BH OF C_60 IS
SIGNAL	clk_out:	STD_LOGIC;
SIGNAL	c1,c0:	STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	c1 <= DIN(7 DOWNTO 4);
	c0 <= DIN(3 DOWNTO 0);
	PROCESS(clk)
	BEGIN
		IF (CLK'EVENT AND clk='1') THEN
			IF (c1=5 AND c0=9) THEN
				clk_out <= '1';
			ELSE CLK_OUT<='0';
			END IF;
		END IF;
	END PROCESS;
	clk_60 <= clk_out;
END BH;