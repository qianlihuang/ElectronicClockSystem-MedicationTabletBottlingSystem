LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DISPLAY_7 IS
	PORT(DIN:IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		DISPLAY_OUT:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END DISPLAY_7;

ARCHITECTURE BH OF DISPLAY_7 IS
BEGIN
	PROCESS(DIN)
	BEGIN
		IF(DIN(3 DOWNTO 0)="0000")THEN
			DISPLAY_OUT<="1111110";
		ELSIF(DIN(3 DOWNTO 0)="0001")THEN
			DISPLAY_OUT<="0110000";
		ELSIF(DIN(3 DOWNTO 0)="0010")THEN
			DISPLAY_OUT<="1101101";
		ELSIF(DIN(3 DOWNTO 0)="0011")THEN
			DISPLAY_OUT<="1111001";
		ELSIF(DIN(3 DOWNTO 0)="0100")THEN
			DISPLAY_OUT<="0110011";
		ELSIF(DIN(3 DOWNTO 0)="0101")THEN
			DISPLAY_OUT<="1011011";
		ELSIF(DIN(3 DOWNTO 0)="0110")THEN
			DISPLAY_OUT<="1011111";
		ELSIF(DIN(3 DOWNTO 0)="0111")THEN
			DISPLAY_OUT<="1110000";
		ELSIF(DIN(3 DOWNTO 0)="1000")THEN
			DISPLAY_OUT<="1111111";
		ELSIF(DIN(3 DOWNTO 0)="1001")THEN
			DISPLAY_OUT<="1111011";
		ELSE
			DISPLAY_OUT<="0000000";
		END IF;
	END PROCESS;
END BH;